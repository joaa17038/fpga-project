/Users/shiju/Documents/FPGA/data/testbench.vhd