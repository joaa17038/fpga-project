/Users/shiju/Documents/FPGA/data/project_1/project_1.srcs/sources_1/new/slidingWindowMaximum.vhd